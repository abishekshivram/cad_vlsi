/*************************************************************************************
CS6230:CAD for VLSI Systems - Final Project
Name: Implementation of a configuralble NoC using Python and bluespec
Team Name: Kilbees
Team Members: Abishekshivram AM (EE18B002)
              Gayatri Ramanathan Ratnam (EE18B006)
              Lloyd K L (CS21M001)
Description: The configurable parameters are defined in this file
Last updated on: 09-Dec-2021
**************************************************************************************/

//This file is meant to be generated by Python script

package Parameters;

//Modify here for changing network address length 
typedef UInt#(16) NetAddressLen;

//Modify here for changing node address length 
typedef UInt#(16) NodeAddressLen;

//For payload parameterisation, change the size here
typedef UInt#(64) PayloadLen;

//A type to represet the clock count
typedef PayloadLen ClockCount;

//3 indicates the no of networks (L1 node count). This value will change based on the network count
Integer l1NodeCount=fromInteger(3);

interface MaxAddressInterface;
    method NodeAddressLen getMaxAddress(NetAddressLen index);
endinterface: MaxAddressInterface

(* synthesize *)
module mkMaxAddress(MaxAddressInterface);
    
    //An array supporitng the core module genrate valid filt addresses
    //NodeAddressLen represents the maximum value each array element can store
    //Each element of the array contains the maximum address possible in that L2 network
    NodeAddressLen maxNodeAddress[l1NodeCount];

    //initialise the max address of each network
    maxNodeAddress[0]=fromInteger(6);
    maxNodeAddress[1]=fromInteger(6);
    maxNodeAddress[2]=fromInteger(6);
    //maxNodeAddress[3]=fromInteger(8);
    //maxNodeAddress[4]=fromInteger(12);

    method NodeAddressLen getMaxAddress(NetAddressLen index);
        return maxNodeAddress[index];
    endmethod: getMaxAddress

endmodule: mkMaxAddress

endpackage: Parameters
