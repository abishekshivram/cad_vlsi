/*************************************************************************************
CS6230:CAD for VLSI Systems - Final Project
Name: Implementation of a configuralble NoC using Python and bluespec
Team Name: Kilbees
Team Members: Abishekshivram AM (EE18B002)
              Gayatri Ramanathan Ratnam (EE18B006)
              Lloyd K L (CS21M001)
Description: Implementation of core - which generates valid flits in random, and consumes flit destined to it
Last updated on: 09-Dec-2021
**************************************************************************************/

package Core;

import Parameters::*;
import Shared::*;
import FIFO::*;
import LFSR::*;

// Interface for the core module 
// Implements methods to get the valid flit generated by the core and to consume the flits destined to this core
interface CoreInterface;

    // A method to check if this core has a valid flit to supply -returns True/False
    method Bool is_flit_generated();

    //Returns the generated flit currently in the core's buffer
    method Flit get_generated_flit();

    // Method to assign a flit to be consumed by this core
    method Action put_flit(Flit flit);

endinterface: CoreInterface

// Implementation of the core module. Mainly implements a rule which generates the flits randomly in different clock cycles.
// Accepts two paraneters - Address of 'this' node and the head node address of the network to which this node (core) belongs
// These two parameters are used to set source address and current destination fields in the generated flit

(* synthesize *)
module mkCore#(parameter Address sourceAddress, parameter Address head_node_addr ) (CoreInterface);

    Reg#(Flit) flitReg          <- mkReg(?); //Uninitialised register to store generated flit
    Reg#(Bool) flitValidStat    <- mkReg(False); //To indicate the content of flitReg is valid or not
    Reg#(Address) myAddress     <- mkReg(sourceAddress); //Register storing the Address of this Core/Node
    Reg#(Address) head_node_address <- mkReg(head_node_addr); //Register storing the Address of this Core/Node

    FIFO#(Flit) flit_consume_fifo   <- mkFIFO; //A fifo to store the consumed flit

    // Set of Lnear Feedback Shift Registers for generating random patterns
    // Used in random rule firing and random destination address generation
    LFSR#(Bit#(16)) lfsr            <- mkLFSR_16; //Helps in firig the flit generation rule randomly
    LFSR#(Bit#(8)) lfsrNodeX        <- mkLFSR_8;  //Helps in generating destination address randomly
    LFSR#(Bit#(8)) lfsrNodeY        <- mkLFSR_8;
    LFSR#(Bit#(8)) lfsrNetX         <- mkLFSR_8;
    LFSR#(Bit#(8)) lfsrNetY         <- mkLFSR_8;
    
    //A flag which helps to fire the fireOnce rule only once.
    // Used to initialise the Lnear Feedback Shift Registers
    Reg#(Bool) fireOnceFlag     <- mkReg(True); 
    Reg#(ClockCount) clockCount <- mkReg(0); //A register to store the clock pulse count
    
    MaxAddressInterface addressLengths <- mkMaxAddress; //instantiates mkMaxAddress from Parameters package


    //A rule to fire only once to seed the different LFSRs
    (* preempts = "fireOnce, (generateFlit,resetFlitStat)" *)
    rule fireOnce (fireOnceFlag);
        fireOnceFlag <= False;
        lfsr.seed('h19);
        lfsrNodeX.seed('h03);
        lfsrNodeY.seed('h11);
        lfsrNetX.seed('h13);
        lfsrNetY.seed('h17);
    endrule

    //Counts the clock pulse, always fire
    rule clockCounter;
        clockCount <= clockCount+1;
        if(myAddress.nodeAddress==fromInteger(0) && myAddress.netAddress==fromInteger(0)) // To prevent all the cores from printing the same statement
            $display("\nClock Cycle: %d",clockCount);
    endrule

    // This rule fires randomly for different core instantiations (32768=(2^16)/2)
    // This is meant for generating valid flits randomly
    (* preempts = "generateFlit, resetFlitStat" *)
    rule generateFlit(lfsr.value() < 32768); 

    //rule generateFlit(clockCount==3 || clockCount==8 || clockCount==11); //NOTE for testing. 
        //if(myAddress.nodeAddress==fromInteger(0) && myAddress.netAddress==fromInteger(0)) //NOTE Test line: Generate flit from Node 0 only.
            //begin
                
                Flit flit;
                flit.srcAddress.netAddress          = myAddress.netAddress;
                flit.srcAddress.nodeAddress         = myAddress.nodeAddress;

                NetAddressX destNetAddressX         = fromInteger(0);
                if(addressLengths.getMaxNetAddressX()!=0) begin //maxNetAddressX,maxNetAddressY can be zero, To handle division by zero
                    destNetAddressX                 = unpack(lfsrNetX.value()%pack(addressLengths.getMaxNetAddressX())); 
                end

                NetAddressY destNetAddressY         = fromInteger(0);
                if(addressLengths.getMaxNetAddressY()!=0) begin 
                    destNetAddressY                 = unpack(lfsrNetY.value()%pack(addressLengths.getMaxNetAddressY())); 
                end

                let destNetAddress                  = {destNetAddressY,destNetAddressX};
                flit.finalDstAddress.netAddress     = destNetAddress;

                NetAddressY l2_array_index = ((addressLengths.getMaxNetAddressX())*destNetAddressY)+destNetAddressX; //NetAddressY type acts just like an int to access aray element

                NodeAddressX destNodeAddressX       = fromInteger(0);
                if(addressLengths.getMaxAddressX(l2_array_index)!=0) begin
                    destNodeAddressX                = unpack(lfsrNodeX.value()%pack(addressLengths.getMaxAddressX(l2_array_index)));
                end
                NodeAddressY destNodeAddressY       = fromInteger(0);
                if(addressLengths.getMaxAddressY(l2_array_index)!=0) begin
                    destNodeAddressY                = unpack(lfsrNodeY.value()%pack(addressLengths.getMaxAddressY(l2_array_index)));
                end
                
                NodeAddress destNodeAddress         = {destNodeAddressY,destNodeAddressX};
                flit.finalDstAddress.nodeAddress    = destNodeAddress;

                if(flit.srcAddress.netAddress==flit.finalDstAddress.netAddress) begin
                    flit.currentDstAddress.netAddress   = flit.finalDstAddress.netAddress;
                    flit.currentDstAddress.nodeAddress  = flit.finalDstAddress.nodeAddress;
                end
                else begin
                    flit.currentDstAddress.netAddress   = head_node_address.netAddress;
                    flit.currentDstAddress.nodeAddress  = head_node_address.nodeAddress;
                end
                
                flit.payload                        = clockCount;

                flitReg                             <= flit;
                if(myAddress!=flit.finalDstAddress) begin //Generate only the flits which are not self destined 
                    flitValidStat                   <= True;
                    $display("Flit generated | Source: %d (Network),%d (Node) | Destination: -> %d (Network),%d (Node)",flit.srcAddress.netAddress,flit.srcAddress.nodeAddress,flit.finalDstAddress.netAddress,flit.finalDstAddress.nodeAddress);
                end    

            //end
        lfsr.next();
        lfsrNodeX.next();
        lfsrNodeY.next();
        lfsrNetX.next();
        lfsrNetY.next();
    endrule

    // If the generateFlit rule is not fired, this rule sets the flit as invalid one
    // Indicating that the flit currently in the 'flitReg' is invalid (Already used)
    rule resetFlitStat;
        flitValidStat <= False;
        lfsr.next();
        lfsrNodeX.next();
        lfsrNodeY.next();
        lfsrNetX.next();
        lfsrNetY.next();
    endrule
    
    // NOTE This rule can add additional delay to other flits which is waiting to be writtten to this fifo (consume fifo)
    // This rule has the highest priority
    // This rule calculates the total flit transmission delay in clock cycle counts
    (* descending_urgency = "calculateDelay" *)
    rule calculateDelay;
        let flit=flit_consume_fifo.first(); flit_consume_fifo.deq();
        $display("############## Transmission Delay: %d, Payload: %d | %d,%d->%d,%d|", clockCount-flit.payload,flit.payload,flit.srcAddress.netAddress,flit.srcAddress.nodeAddress,flit.finalDstAddress.netAddress,flit.finalDstAddress.nodeAddress);
    endrule:calculateDelay

    // Method to check if a valid flit is generated or not
    method Bool is_flit_generated();
        return flitValidStat;
    endmethod

    // Method to get the flit in the flit register
    method Flit get_generated_flit();
        return flitReg;
    endmethod

    // A method to store the flit destined for this core (node)
    method Action put_flit(Flit flit);
        flit_consume_fifo.enq(flit);
        $display(">>>>>>>>>>>>>>> Flit received with payload: %h  | Source: %h (Network),%h (Node) | Destination: -> %h (Network),%h (Node) | MyAddress: -> %h (Network),%h (Node)",          flit.payload,flit.srcAddress.netAddress,flit.srcAddress.nodeAddress,flit.finalDstAddress.netAddress,flit.finalDstAddress.nodeAddress,myAddress.netAddress,myAddress.nodeAddress);
    endmethod

    
endmodule: mkCore

endpackage: Core
