/*************************************************************************************
CS6230:CAD for VLSI Systems - Final Project
Name: Implementation of a configuralble NoC using Python and bluespec
Team Name: Kilbees
Team Members: Abishekshivram AM (EE18B002)
              Gayatri Ramanathan Ratnam (EE18B006)
              Lloyd K L (CS21M001)
Description: The configurable parameters are defined in this file
Last updated on: 09-Dec-2021
**************************************************************************************/

//This file is meant to be generated by Python script

package Parameters;

//Modify here for changing network address length 
typedef Int#(16) NetAddressLen;

//Modify here for changing node address length 
typedef Int#(16) NodeAddressLen;

//For payload parameterisation, change the size here
typedef Int#(16) PayloadLen;

(* synthesize *)
module mkMaxAddress(Empty);
    //An array supporitng the core module genrate valid filt addresses
    //NodeAddressLen represents the maximum value each array element can store
    //5 indicates the no of networks (L1 node count). This value will change based on the network count
    //Each element of the array contains the maximum address possible in that L2 network
    NodeAddressLen maxNodeAddress[5];
    //initialise the max address of each network
    maxNodeAddress[0]=fromInteger(6);
    maxNodeAddress[1]=fromInteger(16);
    maxNodeAddress[2]=fromInteger(4);
    maxNodeAddress[3]=fromInteger(8);
    maxNodeAddress[4]=fromInteger(12);

endmodule: mkMaxAddress

endpackage: Parameters
