/*************************************************************************************
CS6230:CAD for VLSI Systems - Final Project
Name: Implementation of a configuralble NoC using Python and bluespec
Team Name: Kilbees
Team Members: Abishekshivram AM (EE18B002)
              Gayatri Ramanathan Ratnam (EE18B006)
              Lloyd K L (CS21M001)
Description: Represents a node in a chain based network
Last updated on: 09-Dec-2021
**************************************************************************************/

package ChainNodeL2HeadVC;

import Shared::*;
import Parameters::*;

import FIFO :: * ;
import Core :: * ;
import ChainRouterL2HeadVC :: *;


// Interface exposed by the Chain Head Node
// This interface is used by the NoC to build interconnection between nodes
interface IfcChainL2HeadNode;

    // Methods to put flits to the input link buffer of the router. 
    // Each input link has one associated router. Core of the node too has an associated router.
    // Flits that come from left neighbour are inserted to the node's router_left's input link buffer
    // Flits that come from right neighbour are inserted to the node's router_rights's input link buffer
    // Flits that come from L1 neighbour are inserted to the node's L1 input link buffer
    method Action put_value_from_l1(Flit data_from_L1);
    method Action put_value_from_left(Flit data_left);
    method Action put_value_from_right(Flit data_right);

    // Get Value is used to read the value from the respective router
    method ActionValue#(Flit) get_value_to_l1();
    method ActionValue#(Flit) get_value_to_left();
    method ActionValue#(Flit) get_value_to_right();

endinterface


// Module to implement the chain head node.
// This module mainly inplements the rules implementing the round robin arbiter for the output link VCs
// Accepts two parameters - source address and current destination to be used in flit and for flit routing 

(* synthesize *)
module mkChainL2HeadNode #(parameter Address my_addr, parameter Address head_node_addr ) (IfcChainL2HeadNode);


    // Core and four routers - core, left link, right link  and L1 instantiation
    let core            <- mkCore(my_addr,head_node_addr); 
    let router_left     <- mkChainRouterL2HeadVC(my_addr); // takes input from left neighbour and puts in corresponding VC
    let router_right    <- mkChainRouterL2HeadVC(my_addr);
    let router_core     <- mkChainRouterL2HeadVC(my_addr);
    let router_L1       <- mkChainRouterL2HeadVC(my_addr);

    // FIFOs to store the flits from VCs to be moved to the output links present in the node.
    FIFO#(Flit) output_link_left    <- mkFIFO;
    FIFO#(Flit) output_link_right   <- mkFIFO;
    FIFO#(Flit) output_link_l1      <- mkFIFO;

    // This counter is used by arbiters to choose VC to send out data
    // This counter helps to fire different arbiter rules in a round robin fashion 
    Reg#(Bit#(3)) counter   <- mkReg(0);
    rule count_every_cycle;
        if(counter == 3'b101) counter <= 0;
        else counter <= counter + 1;
    endrule

    // Rule to move the valid flit generated by the core to the core-router
    rule core_to_router;
        let flit_generated = core.get_generated_flit();
        if(core.is_flit_generated()==True)
            router_core.put_value(flit_generated);
    endrule

    //A counter to help deciding when to display link utilisation
    // This is a clock interval for printing the link utilisation
    Reg#(LinkUtiliPrInterval) link_util_print_interval <- mkReg(0); 
    rule incr_link_util_print_interval;
        link_util_print_interval <= link_util_print_interval+1;
    endrule

    // This rule prints the link utilisation of the link associated with this node 
    // when the LinkUtiliPrInterval counter is reset
    rule print_link_utilisation(link_util_print_interval==0);
        let rl=router_left.get_link_util_counter();
        let rr=router_right.get_link_util_counter();
        let rl1=router_L1.get_link_util_counter();
        $display("@@@@@@@@@@@@@@@ Link utilisation at Node:%h,%h | : Left Link->%d, Right Link->%d, L1 Link->%d",my_addr.netAddress,my_addr.nodeAddress,rl,rr,rl1);
    endrule
    

    // These six rules are used to move data from router left, L1 router and router rights VCs (VC1 & VC2) to the core router
    // VC1 and VC2 are used to send data to the core 
    // In this rule, we choose VC1 or VC2 from router_left or router_right in a round robin fashion (implemented through 3 bit counter) 
    rule outputLinkCore0(counter == 3'b000);
        $display("here flit is put into core from router left vc1; Arbiter count-%d", counter);      
        Flit data_core=defaultValue;
        data_core <- router_left.get_valueVC1();
        core.put_flit(data_core);
    endrule
    
    rule outputLinkCore1(counter == 3'b001);
        $display("here flit is put into core from router_right vc1; Arbiter count-%d", counter);      
        Flit data_core=defaultValue;
        data_core <- router_right.get_valueVC1();
        core.put_flit(data_core);
    endrule

    rule outputLinkCore2(counter == 3'b010);
        $display("here flit is put into core from router_right vc1; Arbiter count-%d", counter);      
        Flit data_core=defaultValue;
        data_core <- router_L1.get_valueVC1();
        core.put_flit(data_core);
    endrule

    rule outputLinkCore3(counter == 3'b011);
        $display("here flit is put into core from router_left vc2; Arbiter count-%d", counter);      
        Flit data_core=defaultValue;
        data_core <- router_left.get_valueVC2();
        core.put_flit(data_core);
    endrule

    rule outputLinkCore4(counter == 3'b100);
        $display("here flit is put into core from router_right vc2; Arbiter count-%d", counter);      
        Flit data_core=defaultValue;
        data_core <- router_right.get_valueVC2();
        core.put_flit(data_core);
    endrule
    
    rule outputLinkCore5(counter == 3'b101);
        $display("here flit is put into core from router_right vc2; Arbiter count-%d", counter);      
        Flit data_core=defaultValue;
        data_core <- router_L1.get_valueVC2();
        core.put_flit(data_core);
    endrule


    
    // These six rules are used to move data from router left, router L1 and router core's VCs (VC5 & VC6) to the right output link
    // VC5 and VC6 are used to send data to the right output link
    // In this rule, we choose VC5 or VC6 from router_left, router L1 or router_core in a round robin fashion (implemented through 3 bit counter) 
    rule add_to_link_right0(counter == 3'b000);
        $display("add_to_link_right0-> my_addr %d",my_addr.netAddress);    
        Flit data_right=defaultValue;
        data_right <- router_core.get_valueVC5();
        output_link_right.enq(data_right);
    endrule

    rule add_to_link_right1(counter == 3'b001);
        $display("add_to_link_right1-> my_addr %d",my_addr.netAddress);    
        Flit data_right=defaultValue;
        data_right <- router_left.get_valueVC5();
        output_link_right.enq(data_right);
    endrule

    rule add_to_link_right2(counter == 3'b010);
        $display("add_to_link_right1-> my_addr %d",my_addr.netAddress);    
        Flit data_right=defaultValue;
        data_right <- router_L1.get_valueVC5();
        output_link_right.enq(data_right);
    endrule
    
    rule add_to_link_right3(counter == 3'b011);
        $display("add_to_link_right2-> my_addr %d",my_addr.netAddress);    
        Flit data_right=defaultValue;
        data_right <- router_core.get_valueVC6();
        output_link_right.enq(data_right);
    endrule

    rule add_to_link_right4(counter == 3'b100);
        $display("add_to_link_right3-> my_addr %d",my_addr.netAddress);    
        Flit data_right=defaultValue;
        data_right <- router_left.get_valueVC6();
        output_link_right.enq(data_right);
    endrule
    
    rule add_to_link_right5(counter == 3'b101);
        $display("add_to_link_right0-> my_addr %d",my_addr.netAddress);    
        Flit data_right=defaultValue;
        data_right <- router_L1.get_valueVC6();
        output_link_right.enq(data_right);
    endrule


    // These six rules are used to move data from router right, router L1 and router core's VCs (VC3 & VC4) to the left output link
    // VC3 and VC4 are used to send data to the left output link
    // In this rule, we choose VC3 or VC4 from router_right, router L1 or router_core in a round robin fashion (implemented through 3 bit counter) 
    rule add_to_link_left0(counter == 3'b000);
        $display("add_to_link_left0 -> my_addr %d",my_addr.netAddress);    
        Flit data_left=defaultValue;
        data_left <- router_right.get_valueVC3();
        output_link_left.enq(data_left);
    endrule

    rule add_to_link_left1(counter == 3'b001);
        $display("add_to_link_left1 -> my_addr %d",my_addr.netAddress);    
        Flit data_left=defaultValue;
        data_left <- router_core.get_valueVC3();
        output_link_left.enq(data_left);
    endrule

    rule add_to_link_left2(counter == 3'b010);
        $display("add_to_link_left1 -> my_addr %d",my_addr.netAddress);    
        Flit data_left=defaultValue;
        data_left <- router_L1.get_valueVC3();
        output_link_left.enq(data_left);
    endrule
    
    rule add_to_link_left3(counter == 3'b011);
        $display("add_to_link_left2 -> my_addr %d",my_addr.netAddress);    
        Flit data_left=defaultValue;
        data_left <- router_right.get_valueVC4();
        output_link_left.enq(data_left);
    endrule

    rule add_to_link_left4(counter == 3'b100);
        $display("add_to_link_left3 -> my_addr %d",my_addr.netAddress);    
        Flit data_left=defaultValue;
        data_left <- router_core.get_valueVC4();
        output_link_left.enq(data_left);
    endrule

    rule add_to_link_left5(counter == 3'b101);
        $display("add_to_link_left3 -> my_addr %d",my_addr.netAddress);    
        Flit data_left=defaultValue;
        data_left <- router_L1.get_valueVC4();
        output_link_left.enq(data_left);
    endrule


    // These six rules are used to move data from router right, router left and router core's VCs (VC7 & VC8) to the L1 output link
    // VC7 and VC8 are used to send data to the L1 output link
    // In this rule, we choose VC7 or VC7 from router_right, router left or router_core in a round robin fashion (implemented through 3 bit counter) 
    rule add_to_link_l10(counter == 3'b000);
        $display("add_to_link_l10-> my_addr %d",my_addr.netAddress);    
        Flit data_right=defaultValue;
        data_right <- router_core.get_valueVC7();
        output_link_l1.enq(data_right);
    endrule

    rule add_to_link_l11(counter == 3'b001);
        $display("add_to_link_l11-> my_addr %d",my_addr.netAddress);    
        Flit data_right=defaultValue;
        data_right <- router_left.get_valueVC7();
        output_link_l1.enq(data_right);
    endrule

    rule add_to_link_l12(counter == 3'b010);
        $display("add_to_link_l11-> my_addr %d",my_addr.netAddress);    
        Flit data_right=defaultValue;
        data_right <- router_right.get_valueVC7();
        output_link_l1.enq(data_right);
    endrule
    
    rule add_to_link_l13(counter == 3'b011);
        $display("add_to_link_l12-> my_addr %d",my_addr.netAddress);    
        Flit data_right=defaultValue;
        data_right <- router_core.get_valueVC8();
        output_link_l1.enq(data_right);
    endrule

    rule add_to_link_l14(counter == 3'b100);
        $display("add_to_link_l13-> my_addr %d",my_addr.netAddress);    
        Flit data_right=defaultValue;
        data_right <- router_left.get_valueVC8();
        output_link_l1.enq(data_right);
    endrule
    
    rule add_to_link_l15(counter == 3'b101);
        $display("add_to_link_l10-> my_addr %d",my_addr.netAddress);    
        Flit data_right=defaultValue;
        data_right <- router_right.get_valueVC8();
        output_link_l1.enq(data_right);
    endrule

    // Methods to get the flit from output link and return
    // These methods are invoked by the NoC module to make connections between nodes

    // Method to take the flit from left output link and return 
    method ActionValue#(Flit) get_value_to_left();
        let data_to_left = output_link_left.first();
        output_link_left.deq();
        return data_to_left;
    endmethod

    // Method to take the flit from right output link and return 
    method ActionValue#(Flit) get_value_to_right();
        let data_to_right = output_link_right.first();
        output_link_right.deq();
        return data_to_right;
    endmethod

    // Method to take the flit from L1 output link and return 
    method ActionValue#(Flit) get_value_to_l1();
        let data_to_l1 = output_link_l1.first();
        output_link_l1.deq();
        return data_to_l1;
    endmethod

    // Methods to put flits to the input link buffer of the router. 
    // Each input link has one associated router. Core of the node too has an associated router.

    // The flits that come from L1 neighbour are inserted to the node's L1 router input link buffer
    method Action put_value_from_l1(Flit data_from_L1);
        router_L1.put_value(data_from_L1);
    endmethod

    // The flits that come from left neighbour are inserted to the node's router_left's input link buffer
    method Action put_value_from_left(Flit data_left);
        router_left.put_value(data_left);
    endmethod

    // The flits that come from right neighbour are inserted to the router_right's input link buffer
    method Action put_value_from_right(Flit data_right);
        router_right.put_value(data_right);
    endmethod

  
endmodule

endpackage: ChainNodeL2HeadVC
